module special_one_pulse (
    input wire clk,
    input wire pb_in,
    output reg pb_out
);

reg[9:0] pb_in_delay;

always @(posedge clk) begin
	if (pb_in == 1 && pb_in_delay == 0) begin
		pb_out <= 1;
	end 
	else begin
		pb_out <= 0;
	end
end

always @(posedge clk) begin
	pb_in_delay <= {pb_in_delay[8:0] ,pb_in};
end

endmodule

module debounce (
	input wire clk,
	input wire pb, 
	output wire pb_debounced 
);
	reg [3:0] shift_reg; 

	always @(posedge clk) begin
		shift_reg[3:1] <= shift_reg[2:0];
		shift_reg[0] <= pb;
	end

	assign pb_debounced = ((shift_reg == 4'b1111) ? 1'b1 : 1'b0);

endmodule


module one_pulse (
    input wire clk,
    input wire pb_in,
    output reg pb_out
);

	reg pb_in_delay;

	always @(posedge clk) begin
		if (pb_in == 1'b1 && pb_in_delay == 1'b0) begin
			pb_out <= 1'b1;
		end else begin
			pb_out <= 1'b0;
		end
	end
	
	always @(posedge clk) begin
		pb_in_delay <= pb_in;
	end
endmodule
